package UMDRISC_PKG is

	CONSTANT DATA_WIDTH:INTEGER := 24;
	CONSTANT ADDRESS_WIDTH:INTEGER := 24;
	CONSTANT PC_WIDTH:INTEGER := 24;

end UMDRISC_PKG;

package body UMDRISC_PKG is

end UMDRISC_PKG;
