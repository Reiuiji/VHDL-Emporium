------------------------------------------------------------
-- implemented the 8 Byte X 24 byte memory
--
-- Instruction memory on it is the following:
--
-- ADDI  R0, 2   ; ADDI R0<-2           500002
-- ADDI  R1, 1   ; ADDI R1<-1           510001
-- ADD   R0, R1  ; ADD  R0<-R0 + R1     001000
-- AND   R0, R1  ; AND  R0<-R0 & R1     201000
-- OR    R0, R1  ; OR   R0<-R0 or R1    301000
-- ADD   R0, R1  ; ADD  R0<-R0 + R1     001000
-- MOV   R5, R0  ; R5 <- R0             450000
--
-----------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity RAM_8x24 is
	generic(
		RAM_WIDTH:	integer:=8; -- 00 - FF choice
		DATA_WIDTH: integer:=24
	);
	port(
		CLOCK			: in std_logic;
		WE				: in std_logic;
        --OUTPUT RAM
		OUT_ADDR		: in std_logic_vector(RAM_WIDTH-1 downto 0);
		OUT_DATA		: out std_logic_vector(DATA_WIDTH-1 downto 0);
		--INPUT RAM
		IN_ADDR		    : in std_logic_vector(RAM_WIDTH-1 downto 0);
		IN_DATA			: in std_logic_vector(DATA_WIDTH-1 downto 0)
   );
end RAM_8x24;

architecture RAM_ARCH of RAM_8x24 is

	type    ram_type is array (0 to 2**RAM_WIDTH-1) of std_logic_vector (DATA_WIDTH-1 downto 0);
    signal  RAM : ram_type := (
		x"500002", x"510001", x"001000", x"201000", x"301000", x"001000", x"450000", x"000000", -- 00 - 07
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- 08 - 0F
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- 10 - 17
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- 18 - 1F
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- 20 - 27
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- 28 - 2F
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- 30 - 37
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- 38 - 3F
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- 40 - 47
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- 48 - 4F
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- 50 - 57
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- 58 - 5F
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- 60 - 67
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- 68 - 6F
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- 70 - 77
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- 78 - 7F
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- 80 - 87
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- 88 - 8F
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- 90 - 97
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- 98 - 9F
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- A0 - A7
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- A8 - AF
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- B0 - B7
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- B8 - BF
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- C0 - C7
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- C8 - CF
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- D0 - D7
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- D8 - DF
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- E0 - E7
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- E8 - EF
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", -- F0 - F7
		x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000", x"000000"  -- F8 - FF
	);


	signal	ADDR_IN: std_logic_vector(RAM_WIDTH-1 downto 0);
	
begin
   process(CLOCK,WE)
   begin
			if (CLOCK'event and CLOCK = '0') then
				if (WE = '1') then
					RAM(to_integer(unsigned(IN_ADDR))) <= IN_DATA;
				end if;
				ADDR_IN <= OUT_ADDR;
			end if;
	end process;
	OUT_DATA <= RAM(to_integer(unsigned(ADDR_IN)));
end RAM_ARCH;
